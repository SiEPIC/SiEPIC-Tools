* Spice output from KLayout SiEPIC-Tools v0.3.12, 2018-01-21 12:18:56.

.subckt GSiP_RingMod_Transceiver Ring_Modulator_DB_1_elec1a Ring_Modulator_DB_1_elec1c Ring_Modulator_DB_1_elec2h1 Ring_Modulator_DB_1_elec2h2 Ring_Modulator_DB_2_elec1a Ring_Modulator_DB_2_elec1c Ring_Modulator_DB_2_elec2h1 Ring_Modulator_DB_2_elec2h2 Ring_Modulator_DB_3_elec1a Ring_Modulator_DB_3_elec1c Ring_Modulator_DB_3_elec2h1 Ring_Modulator_DB_3_elec2h2 Ring_Modulator_DB_4_elec1a Ring_Modulator_DB_4_elec1c Ring_Modulator_DB_4_elec2h1 Ring_Modulator_DB_4_elec2h2 Detector_Ge_floating_4_elecN Detector_Ge_floating_4_elecP Detector_Ge_floating_5_elecN Detector_Ge_floating_5_elecP Detector_Ge_floating_6_elecN Detector_Ge_floating_6_elecP Detector_Ge_floating_7_elecN Detector_Ge_floating_7_elecP Ring_Filter_DB_3_elec2h1 Ring_Filter_DB_3_elec2h2 Ring_Filter_DB_4_elec2h1 Ring_Filter_DB_4_elec2h2 Ring_Filter_DB_2_elec2h1 Ring_Filter_DB_2_elec2h2 Ring_Filter_DB_1_elec2h1 Ring_Filter_DB_1_elec2h2 Detector_Ge_floating_27_elecN Detector_Ge_floating_27_elecP Detector_Ge_floating_28_elecN Detector_Ge_floating_28_elecP Detector_Ge_floating_29_elecN Detector_Ge_floating_29_elecP Detector_Ge_floating_30_elecN Detector_Ge_floating_30_elecP edgecoupler_1550_laser1 edgecoupler_1550_detector3 edgecoupler_1550_detector2
.param MC_uniformity_width=0 
.param MC_uniformity_thickness=0 
.param MC_resolution_x=100 
.param MC_resolution_y=100 
.param MC_grid=10e-6 
.param MC_non_uniform=99 
 Ring_Modulator_DB_1  Ring_Modulator_DB_1_elec1a Ring_Modulator_DB_1_elec1c Ring_Modulator_DB_1_elec2h1 Ring_Modulator_DB_1_elec2h2 N$3 N$2 N$1 N$0 Ring_Modulator_DB library="Design kits/GSiP" radius=10.000u wg_width=0.500u gap=0.310u gap_monitor=0.450u lay_x=2.14E-3 lay_y=612.175E-6 sch_x=13.917513641E0 sch_y=3.981286875E0 
 Ring_Modulator_DB_2  Ring_Modulator_DB_2_elec1a Ring_Modulator_DB_2_elec1c Ring_Modulator_DB_2_elec2h1 Ring_Modulator_DB_2_elec2h2 N$6 N$7 N$5 N$4 Ring_Modulator_DB library="Design kits/GSiP" radius=10.025u wg_width=0.500u gap=0.310u gap_monitor=0.450u lay_x=2.59E-3 lay_y=612.2E-6 sch_x=16.844093612E0 sch_y=3.981449463E0 
 Ring_Modulator_DB_3  Ring_Modulator_DB_3_elec1a Ring_Modulator_DB_3_elec1c Ring_Modulator_DB_3_elec2h1 Ring_Modulator_DB_3_elec2h2 N$11 N$8 N$10 N$9 Ring_Modulator_DB library="Design kits/GSiP" radius=10.050u wg_width=0.500u gap=0.310u gap_monitor=0.450u lay_x=3.04E-3 lay_y=612.225E-6 sch_x=19.770673583E0 sch_y=3.981612051E0 
 Ring_Modulator_DB_4  Ring_Modulator_DB_4_elec1a Ring_Modulator_DB_4_elec1c Ring_Modulator_DB_4_elec2h1 Ring_Modulator_DB_4_elec2h2 N$12 N$15 N$14 N$13 Ring_Modulator_DB library="Design kits/GSiP" radius=10.075u wg_width=0.500u gap=0.310u gap_monitor=0.450u lay_x=3.49E-3 lay_y=612.25E-6 sch_x=22.697253554E0 sch_y=3.981774639E0 
 Detector_Ge_floating_4  Detector_Ge_floating_4_elecN Detector_Ge_floating_4_elecP N$16 Detector_Ge_floating library="Design kits/GSiP"  lay_x=150.0E-6 lay_y=585.95E-6 sch_x=975.526657E-3 sch_y=3.810732298E0  sch_r=90
 Detector_Ge_floating_5  Detector_Ge_floating_5_elecN Detector_Ge_floating_5_elecP N$17 Detector_Ge_floating library="Design kits/GSiP"  lay_x=250.0E-6 lay_y=525.95E-6 sch_x=1.625877762E0 sch_y=3.420521635E0  sch_r=90
 Detector_Ge_floating_6  Detector_Ge_floating_6_elecN Detector_Ge_floating_6_elecP N$18 Detector_Ge_floating library="Design kits/GSiP"  lay_x=350.0E-6 lay_y=465.95E-6 sch_x=2.276228866E0 sch_y=3.030310972E0  sch_r=90
 Detector_Ge_floating_7  Detector_Ge_floating_7_elecN Detector_Ge_floating_7_elecP N$19 Detector_Ge_floating library="Design kits/GSiP"  lay_x=450.0E-6 lay_y=405.95E-6 sch_x=2.926579971E0 sch_y=2.64010031E0  sch_r=90
 wg_strip_integral_1550_8  N$8 N$12 wg_strip_integral_1550 library="Design kits/GSiP" wg_length=405.375u wg_width=0.500u points=[[3062.3,820.52],[3467.675,820.52]] radius=5.0 lay_x=3.264987E-3 lay_y=600.52E-6 sch_x=21.233879023E0 sch_y=3.905488454E0 
 terminator_te1550_9  N$0 terminator_te1550 library="Design kits/GSiP"  lay_x=2.1677E-3 lay_y=622.28E-6 sch_x=14.097660897E0 sch_y=4.047004854E0  sch_r=180
 terminator_te1550_10  N$4 terminator_te1550 library="Design kits/GSiP"  lay_x=2.617725E-3 lay_y=622.33E-6 sch_x=17.024403456E0 sch_y=4.04733003E0  sch_r=180
 terminator_te1550_11  N$9 terminator_te1550 library="Design kits/GSiP"  lay_x=3.06775E-3 lay_y=622.38E-6 sch_x=19.951146015E0 sch_y=4.047655206E0  sch_r=180
 terminator_te1550_12  N$13 terminator_te1550 library="Design kits/GSiP"  lay_x=3.517775E-3 lay_y=622.43E-6 sch_x=22.877888574E0 sch_y=4.047980381E0  sch_r=180
 wg_strip_integral_1550_13  N$14 N$16 wg_strip_integral_1550 library="Design kits/GSiP" wg_length=3380.990u wg_width=0.500u points=[[3467.675,842.43],[3261.08,842.43],[3261.08,870.0],[1530.8,870.0],[1530.8,896.44],[150.0,896.44],[150.0,876.4]] radius=5.0 lay_x=1.808212E-3 lay_y=649.435E-6 sch_x=11.759726718E0 sch_y=4.223607697E0 
 wg_strip_integral_1550_14  N$10 N$17 wg_strip_integral_1550 library="Design kits/GSiP" wg_length=2832.479u wg_width=0.500u points=[[3017.7,842.38],[2813.72,842.38],[2813.72,865.0],[250.0,865.0],[250.0,816.4]] radius=5.0 lay_x=1.633225E-3 lay_y=621.325E-6 sch_x=10.62169683E0 sch_y=4.040794001E0 
 wg_strip_integral_1550_15  N$5 N$18 wg_strip_integral_1550 library="Design kits/GSiP" wg_length=2332.554u wg_width=0.500u points=[[2567.725,842.33],[2364.07,842.33],[2364.07,860.0],[350.0,860.0],[350.0,756.4]] radius=5.0 lay_x=1.458237E-3 lay_y=588.825E-6 sch_x=9.483660439E0 sch_y=3.829429892E0 
 wg_strip_integral_1550_16  N$1 N$19 wg_strip_integral_1550 library="Design kits/GSiP" wg_length=1811.483u wg_width=0.500u points=[[2117.75,842.28],[450.0,842.28],[450.0,696.4]] radius=5.0 lay_x=1.28325E-3 lay_y=549.965E-6 sch_x=8.345630551E0 sch_y=3.576703453E0 
 wg_strip_integral_1550_17  N$2 N$6 wg_strip_integral_1550 library="Design kits/GSiP" wg_length=405.475u wg_width=0.500u points=[[2162.25,820.52],[2567.725,820.52]] radius=5.0 lay_x=2.364987E-3 lay_y=600.52E-6 sch_x=15.380719081E0 sch_y=3.905488454E0 
 wg_strip_integral_1550_18  N$7 N$11 wg_strip_integral_1550 library="Design kits/GSiP" wg_length=405.425u wg_width=0.500u points=[[2612.275,820.52],[3017.7,820.52]] radius=5.0 lay_x=2.814987E-3 lay_y=600.52E-6 sch_x=18.307299052E0 sch_y=3.905488454E0 
 terminator_te1550_19  N$34 terminator_te1550 library="Design kits/GSiP"  lay_x=7.58387E-3 lay_y=395.21E-6 sch_x=49.321782325E0 sch_y=2.570252601E0 
 terminator_te1550_20  N$30 terminator_te1550 library="Design kits/GSiP"  lay_x=7.13452E-3 lay_y=395.26E-6 sch_x=46.399429636E0 sch_y=2.570577776E0 
 Ring_Filter_DB_3  Ring_Filter_DB_3_elec2h1 Ring_Filter_DB_3_elec2h2 N$25 N$24 N$22 N$23 Ring_Filter_DB library="Design kits/GSiP" radius=10.050u wg_width=0.500u gap=0.300u gap_monitor=0.320u lay_x=6.71294E-3 lay_y=385.29E-6 sch_x=43.657679449E0 sch_y=2.505737771E0 
 Ring_Filter_DB_4  Ring_Filter_DB_4_elec2h1 Ring_Filter_DB_4_elec2h2 N$29 N$28 N$26 N$27 Ring_Filter_DB library="Design kits/GSiP" radius=10.075u wg_width=0.500u gap=0.300u gap_monitor=0.320u lay_x=6.263595E-3 lay_y=385.315E-6 sch_x=40.735359277E0 sch_y=2.505900359E0 
 terminator_te1550_23  N$22 terminator_te1550 library="Design kits/GSiP"  lay_x=6.68519E-3 lay_y=395.31E-6 sch_x=43.477207017E0 sch_y=2.570902952E0 
 terminator_te1550_24  N$26 terminator_te1550 library="Design kits/GSiP"  lay_x=6.23582E-3 lay_y=395.36E-6 sch_x=40.554724258E0 sch_y=2.571228128E0 
 Ring_Filter_DB_2  Ring_Filter_DB_2_elec2h1 Ring_Filter_DB_2_elec2h2 N$33 N$31 N$30 N$32 Ring_Filter_DB library="Design kits/GSiP" radius=10.025u wg_width=0.500u gap=0.300u gap_monitor=0.320u lay_x=7.162245E-3 lay_y=385.265E-6 sch_x=46.57973948E0 sch_y=2.505575184E0 
 Ring_Filter_DB_1  Ring_Filter_DB_1_elec2h1 Ring_Filter_DB_1_elec2h2 N$35 N$37 N$34 N$36 Ring_Filter_DB library="Design kits/GSiP" radius=10.000u wg_width=0.500u gap=0.300u gap_monitor=0.320u lay_x=7.61157E-3 lay_y=385.24E-6 sch_x=49.501929581E0 sch_y=2.505412596E0 
 Detector_Ge_floating_27  Detector_Ge_floating_27_elecN Detector_Ge_floating_27_elecP N$38 Detector_Ge_floating library="Design kits/GSiP"  lay_x=7.60045E-3 lay_y=617.75E-6 sch_x=49.429610538E0 sch_y=4.017543949E0  sch_r=180
 Detector_Ge_floating_28  Detector_Ge_floating_28_elecN Detector_Ge_floating_28_elecP N$39 Detector_Ge_floating library="Design kits/GSiP"  lay_x=7.15045E-3 lay_y=617.75E-6 sch_x=46.503030567E0 sch_y=4.017543949E0  sch_r=180
 Detector_Ge_floating_29  Detector_Ge_floating_29_elecN Detector_Ge_floating_29_elecP N$40 Detector_Ge_floating library="Design kits/GSiP"  lay_x=6.70045E-3 lay_y=617.75E-6 sch_x=43.576450596E0 sch_y=4.017543949E0  sch_r=180
 Detector_Ge_floating_30  Detector_Ge_floating_30_elecN Detector_Ge_floating_30_elecP N$41 Detector_Ge_floating library="Design kits/GSiP"  lay_x=6.25045E-3 lay_y=617.75E-6 sch_x=40.649870624E0 sch_y=4.017543949E0  sch_r=180
 wg_strip_integral_1550_31  N$35 N$31 wg_strip_integral_1550 library="Design kits/GSiP" wg_length=404.800u wg_width=0.500u points=[[470.68,56.41],[875.48,56.41]] radius=5.0 lay_x=7.38692E-3 lay_y=373.59E-6 sch_x=48.040915824E0 sch_y=2.429646692E0  sch_r=180
 wg_strip_integral_1550_32  N$36 N$38 wg_strip_integral_1550 library="Design kits/GSiP" wg_length=355.526u wg_width=0.500u points=[[426.18,34.79],[339.0,34.79],[339.0,-187.75],[389.1,-187.75]] radius=5.0 lay_x=7.678035E-3 lay_y=506.48E-6 sch_x=49.934185443E0 sch_y=3.293898275E0  sch_r=180
 wg_strip_integral_1550_33  N$32 N$39 wg_strip_integral_1550 library="Design kits/GSiP" wg_length=354.776u wg_width=0.500u points=[[875.48,34.74],[789.0,34.74],[789.0,-187.75],[839.1,-187.75]] radius=5.0 lay_x=7.228385E-3 lay_y=506.505E-6 sch_x=47.0098817E0 sch_y=3.294060863E0  sch_r=180
 wg_strip_integral_1550_34  N$23 N$40 wg_strip_integral_1550 library="Design kits/GSiP" wg_length=354.006u wg_width=0.500u points=[[1324.76,34.69],[1239.0,34.69],[1239.0,-187.75],[1289.1,-187.75]] radius=5.0 lay_x=6.778745E-3 lay_y=506.53E-6 sch_x=44.085642993E0 sch_y=3.294223451E0  sch_r=180
 wg_strip_integral_1550_35  N$27 N$41 wg_strip_integral_1550 library="Design kits/GSiP" wg_length=371.296u wg_width=0.500u points=[[1774.08,34.64],[1679.99,34.64],[1679.99,-187.75],[1739.1,-187.75]] radius=5.0 lay_x=6.33359E-3 lay_y=506.555E-6 sch_x=41.190572533E0 sch_y=3.294386038E0  sch_r=180
 wg_strip_integral_1550_36  N$33 N$24 wg_strip_integral_1550 library="Design kits/GSiP" wg_length=404.730u wg_width=0.500u points=[[920.03,56.41],[1324.76,56.41]] radius=5.0 lay_x=6.937605E-3 lay_y=373.59E-6 sch_x=45.118790758E0 sch_y=2.429646692E0  sch_r=180
 wg_strip_integral_1550_37  N$25 N$28 wg_strip_integral_1550 library="Design kits/GSiP" wg_length=404.720u wg_width=0.500u points=[[1369.36,56.41],[1774.08,56.41]] radius=5.0 lay_x=6.48828E-3 lay_y=373.59E-6 sch_x=42.196600657E0 sch_y=2.429646692E0  sch_r=180
 wg_strip_integral_1550_38  N$3 N$42 wg_strip_integral_1550 library="Design kits/GSiP" wg_length=2413.976u wg_width=0.500u points=[[2117.75,600.52],[1433.8,600.52],[1433.8,100.0],[200.0,100.0]] radius=5.0 lay_x=1.158875E-3 lay_y=350.26E-6 sch_x=7.536756365E0 sch_y=2.277919779E0 
 YBranch_te1550_39  N$43 N$44 N$45 YBranch_te1550 library="Design kits/GSiP"  lay_x=7.415E-3 lay_y=172.0E-6 sch_x=48.223534414E0 sch_y=1.1186039E0 
 edgecoupler_1550_40  edgecoupler_1550_laser1 N$42 edgecoupler_1550 library="Design kits/GSiP"  lay_x=100.0E-6 lay_y=100.0E-6 sch_x=650.351105E-3 sch_y=650.351105E-3 
 edgecoupler_1550_41  edgecoupler_1550_detector3 N$46 edgecoupler_1550 library="Design kits/GSiP"  lay_x=7.75E-3 lay_y=90.0E-6 sch_x=50.402210615E0 sch_y=585.315994E-3  sch_r=180
 edgecoupler_1550_42  edgecoupler_1550_detector2 N$47 edgecoupler_1550 library="Design kits/GSiP"  lay_x=7.75E-3 lay_y=865.0E-6 sch_x=50.402210615E0 sch_y=5.625537056E0  sch_r=180
 wg_strip_integral_1550_43  N$15 N$43 wg_strip_integral_1550 library="Design kits/GSiP" wg_length=4319.401u wg_width=0.500u points=[[3512.325,600.52],[3586.0,600.52],[3586.0,172.0],[7407.5,172.0]] radius=5.0 lay_x=5.459912E-3 lay_y=386.26E-6 sch_x=35.508598008E0 sch_y=2.512046177E0 
 wg_strip_integral_1550_44  N$29 N$47 wg_strip_integral_1550 library="Design kits/GSiP" wg_length=2334.386u wg_width=0.500u points=[[6241.27,373.59],[6022.0,373.59],[6022.0,865.0],[7650.0,865.0]] radius=5.0 lay_x=6.835375E-3 lay_y=619.295E-6 sch_x=44.453936824E0 sch_y=4.027591874E0 
 wg_strip_integral_1550_45  N$44 N$37 wg_strip_integral_1550 library="Design kits/GSiP" wg_length=578.226u wg_width=0.500u points=[[7422.5,174.75],[7720.0,174.75],[7720.0,373.59],[7633.82,373.59]] radius=5.0 lay_x=7.571875E-3 lay_y=274.17E-6 sch_x=49.24377271E0 sch_y=1.783067624E0 
 wg_strip_integral_1550_46  N$45 N$46 wg_strip_integral_1550 library="Design kits/GSiP" wg_length=302.456u wg_width=0.500u points=[[7422.5,169.25],[7582.0,169.25],[7582.0,90.0],[7650.0,90.0]] radius=5.0 lay_x=7.53625E-3 lay_y=129.625E-6 sch_x=49.012085129E0 sch_y=843.017619E-3 
.ends GSiP_RingMod_Transceiver

